// list all paths to your design files
`include "../01_RTL/core.v"
`include "../01_RTL/median_unit.v"
`include "../01_RTL/processing_unit.v"